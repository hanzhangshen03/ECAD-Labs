
module unsaved (
	clk_clk,
	reset_reset_n,
	eightbitstosevenseg_0_led_pins_led0,
	eightbitstosevenseg_0_led_pins_led1);	

	input		clk_clk;
	input		reset_reset_n;
	output	[6:0]	eightbitstosevenseg_0_led_pins_led0;
	output	[6:0]	eightbitstosevenseg_0_led_pins_led1;
endmodule
